

.SUBCKT COMP VCMP_OUT VSTORE VRAMP VDD VSS X1 X2 X3  X4 
MN1 VSS X1 X1 X1 pmos L=1u W=1u
MN2 VSS X1 X2 X2 pmos L=1u W=1u
MN3 X1 VSTORE X3 X3 nmos L=1u W=1u
MN4 X2 VRAMP X3 X3 nmos L=1u W=1u
MN5 X3 V2B VSS VSS nmos L=1u W=1u
MN6 X4 V2B VSS VSS nmos L=1u W=1u
MN7 VSS X2 X4 X4 pmos L=1u W=1u
MN8 VSS X4 VCMP_OUT VCMP_OUT pmos L=1u W=1u
MN9 VCMP_OUT X4 VSS VSS nmos L=1u W=1u
.ENDS