* Comparator testbench
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130_ngspice.spi
.include ../../lib/SUN_TR_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-8 abstol=1e-8

*----------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------

.param TRF = 10n
.param TCLK = 100n
.param C_ERASE = 5
.param C_EXPOSE = 255
.param C_CONVERT = 255
.param C_READ = 5

*- Pulse Width of control signals
.param PW_ERASE =  {(C_ERASE +1)*TCLK}
.param PW_EXPOSE =  {(C_EXPOSE +1)*TCLK}
.param PW_CONVERT =  {(C_CONVERT +1)*TCLK}
.param PW_READ =  {(C_READ +1)*TCLK}

*- Delay of control signals
.param TD_ERASE = {TCLK }
.param TD_EXPOSE = {TD_ERASE + PW_ERASE + TCLK}
.param TD_CONVERT = {TD_EXPOSE + PW_EXPOSE + TCLK}
.param TD_READ = {TD_CONVERT + PW_CONVERT + TCLK}
.param PERIOD = {TD_READ + PW_READ + TCLK}

*- Analog parameters
.param VDD = 1.5
.param VADC_MIN = 0.5
.param VADC_MAX = 1.1
.param VADC_REF = {VADC_MAX - VADC_MIN}
.param VADC_LSB = {VADC_REF/256}

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc VDD
VSS VSS 0 dc 0

*- Control signals
VERASE ERASE 0 dc 0 pulse (0 VDD TD_ERASE TRF TRF PW_ERASE PERIOD)
VEXPOSE EXPOSE 0 dc 0 pulse (0 VDD TD_EXPOSE TRF TRF PW_EXPOSE PERIOD)
VCONVERT CONVERT 0 dc 0 pulse (0 VDD TD_CONVERT TRF TRF PW_CONVERT PERIOD)
VREAD READ 0 dc 0 pulse (0 VDD TD_READ TRF TRF PW_READ PERIOD)

*- ADC related sources
VREF VREF 0 DC VADC_REF
VMAX VMAX 0 DC VADC_MAX
VRESET VRESET VMAX DC 0
VMIN VMIN 0 DC VADC_MIN


*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include comparator.cir

I3 0 VBN1 dc 8u

mnb1 VBN1 VBN1 VSS VSS nmos w=0.5u l=0.5u

VSTORE VSTORE 0 dc 1
XDUT VCMP_OUT VSTORE VRAMP VDD VSS COMP

*----------------------------------------------------------------
* RAMP
*----------------------------------------------------------------
* Use a capacitor and current source to model a ramp
* I = C x dV/dt, where
* dt = PW_CONVERT
* C = 1n
* dV = VADC_MAX - VADC_MIN
BR1 0 VRAMP I = V(CONVERT)*( 1n*(VADC_MAX - VADC_MIN)/PW_CONVERT)
CR1 VRAMP 0 1n ic=0

* SPICE freaks out if any node only have current sources and capacitors on it. so insert a resistor to ground
R1 VRAMP 0 1T

* Model reset as a variable resistor to
BR2 VRAMP VMIN I=V(ERASE)*V(VRAMP,VMIN)/100

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set color0=white
set color1=black
unset askquit
tran 1n 60u
plot V(VRAMP) V(CONVERT) V(ERASE) V(VCMP_OUT)

.endc
.end